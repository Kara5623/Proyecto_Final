module AND(
	input A,B,
	output S
);

assign S= A & B;
endmodule